VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_tx
  CLASS BLOCK ;
  FOREIGN uart_tx ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.385 10.640 26.985 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.115 10.640 61.715 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.845 10.640 96.445 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.575 10.640 131.175 138.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.360 144.680 30.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 61.320 144.680 62.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 93.280 144.680 94.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 125.240 144.680 126.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.060 144.680 27.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 58.020 144.680 59.620 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 89.980 144.680 91.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 121.940 144.680 123.540 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 150.000 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.840 150.000 126.440 ;
    END
  END data_in[7]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END rst_n
  PIN tx_busy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END tx_busy
  PIN tx_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END tx_out
  PIN tx_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 30.640 150.000 31.240 ;
    END
  END tx_start
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 0.070 10.640 144.440 138.960 ;
      LAYER met2 ;
        RECT 0.100 145.720 35.230 146.610 ;
        RECT 36.070 145.720 80.310 146.610 ;
        RECT 81.150 145.720 125.390 146.610 ;
        RECT 126.230 145.720 142.970 146.610 ;
        RECT 0.100 4.280 142.970 145.720 ;
        RECT 0.650 4.000 44.890 4.280 ;
        RECT 45.730 4.000 89.970 4.280 ;
        RECT 90.810 4.000 135.050 4.280 ;
        RECT 135.890 4.000 142.970 4.280 ;
      LAYER met3 ;
        RECT 4.400 139.040 146.000 139.890 ;
        RECT 3.990 126.840 146.000 139.040 ;
        RECT 3.990 125.440 145.600 126.840 ;
        RECT 3.990 92.840 146.000 125.440 ;
        RECT 4.400 91.440 146.000 92.840 ;
        RECT 3.990 79.240 146.000 91.440 ;
        RECT 3.990 77.840 145.600 79.240 ;
        RECT 3.990 45.240 146.000 77.840 ;
        RECT 4.400 43.840 146.000 45.240 ;
        RECT 3.990 31.640 146.000 43.840 ;
        RECT 3.990 30.240 145.600 31.640 ;
        RECT 3.990 10.715 146.000 30.240 ;
      LAYER met4 ;
        RECT 124.495 40.975 124.825 78.705 ;
  END
END uart_tx
END LIBRARY

