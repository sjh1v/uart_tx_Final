module uart_tx (clk,
    rst_n,
    tx_busy,
    tx_out,
    tx_start,
    data_in);
 input clk;
 input rst_n;
 output tx_busy;
 output tx_out;
 input tx_start;
 input [7:0] data_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire \bit_idx[0] ;
 wire \bit_idx[1] ;
 wire \bit_idx[2] ;
 wire \clk_cnt[0] ;
 wire \clk_cnt[10] ;
 wire \clk_cnt[11] ;
 wire \clk_cnt[12] ;
 wire \clk_cnt[13] ;
 wire \clk_cnt[14] ;
 wire \clk_cnt[15] ;
 wire \clk_cnt[1] ;
 wire \clk_cnt[2] ;
 wire \clk_cnt[3] ;
 wire \clk_cnt[4] ;
 wire \clk_cnt[5] ;
 wire \clk_cnt[6] ;
 wire \clk_cnt[7] ;
 wire \clk_cnt[8] ;
 wire \clk_cnt[9] ;
 wire \data_reg[0] ;
 wire \data_reg[1] ;
 wire \data_reg[2] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire parity_bit;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;

 sky130_fd_sc_hd__xnor2_1 _112_ (.A(net2),
    .B(net1),
    .Y(_091_));
 sky130_fd_sc_hd__xnor2_1 _113_ (.A(net8),
    .B(net7),
    .Y(_092_));
 sky130_fd_sc_hd__xnor2_1 _114_ (.A(_091_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__xor2_1 _115_ (.A(net6),
    .B(net5),
    .X(_094_));
 sky130_fd_sc_hd__xnor2_1 _116_ (.A(net4),
    .B(net3),
    .Y(_095_));
 sky130_fd_sc_hd__xnor2_1 _117_ (.A(_094_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_1 _118_ (.A(_093_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__buf_2 _119_ (.A(\state[1] ),
    .X(_098_));
 sky130_fd_sc_hd__nor3_2 _120_ (.A(\state[2] ),
    .B(\state[0] ),
    .C(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__nand2_4 _121_ (.A(net10),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(_097_),
    .A1(net40),
    .S(_100_),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(_101_),
    .X(_000_));
 sky130_fd_sc_hd__inv_2 _124_ (.A(\state[2] ),
    .Y(_102_));
 sky130_fd_sc_hd__mux4_1 _125_ (.A0(\data_reg[0] ),
    .A1(\data_reg[1] ),
    .A2(\data_reg[2] ),
    .A3(\data_reg[3] ),
    .S0(\bit_idx[0] ),
    .S1(\bit_idx[1] ),
    .X(_103_));
 sky130_fd_sc_hd__or2_1 _126_ (.A(\bit_idx[2] ),
    .B(_103_),
    .X(_104_));
 sky130_fd_sc_hd__mux4_1 _127_ (.A0(\data_reg[4] ),
    .A1(\data_reg[5] ),
    .A2(\data_reg[6] ),
    .A3(\data_reg[7] ),
    .S0(\bit_idx[0] ),
    .S1(\bit_idx[1] ),
    .X(_105_));
 sky130_fd_sc_hd__or2b_1 _128_ (.A(_105_),
    .B_N(\bit_idx[2] ),
    .X(_106_));
 sky130_fd_sc_hd__nor2_2 _129_ (.A(\state[2] ),
    .B(\state[0] ),
    .Y(_107_));
 sky130_fd_sc_hd__and2_1 _130_ (.A(_102_),
    .B(\state[0] ),
    .X(_108_));
 sky130_fd_sc_hd__a32o_1 _131_ (.A1(_104_),
    .A2(_106_),
    .A3(_107_),
    .B1(_108_),
    .B2(parity_bit),
    .X(_109_));
 sky130_fd_sc_hd__a2bb2o_1 _132_ (.A1_N(\state[0] ),
    .A2_N(_098_),
    .B1(net12),
    .B2(\state[2] ),
    .X(_110_));
 sky130_fd_sc_hd__a31o_1 _133_ (.A1(_102_),
    .A2(_098_),
    .A3(_109_),
    .B1(_110_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _134_ (.A0(net11),
    .A1(net10),
    .S(_099_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(_111_),
    .X(_002_));
 sky130_fd_sc_hd__or4_1 _136_ (.A(\clk_cnt[3] ),
    .B(\clk_cnt[1] ),
    .C(\clk_cnt[2] ),
    .D(\clk_cnt[0] ),
    .X(_033_));
 sky130_fd_sc_hd__a31o_1 _137_ (.A1(\clk_cnt[5] ),
    .A2(\clk_cnt[4] ),
    .A3(_033_),
    .B1(\clk_cnt[6] ),
    .X(_034_));
 sky130_fd_sc_hd__or4_1 _138_ (.A(\clk_cnt[13] ),
    .B(\clk_cnt[14] ),
    .C(\clk_cnt[12] ),
    .D(\clk_cnt[11] ),
    .X(_035_));
 sky130_fd_sc_hd__or4_1 _139_ (.A(\clk_cnt[10] ),
    .B(\clk_cnt[9] ),
    .C(\clk_cnt[15] ),
    .D(_035_),
    .X(_036_));
 sky130_fd_sc_hd__o21a_1 _140_ (.A1(\state[0] ),
    .A2(\state[1] ),
    .B1(\state[2] ),
    .X(_037_));
 sky130_fd_sc_hd__or2_1 _141_ (.A(_099_),
    .B(_037_),
    .X(_038_));
 sky130_fd_sc_hd__a311o_1 _142_ (.A1(\clk_cnt[8] ),
    .A2(\clk_cnt[7] ),
    .A3(_034_),
    .B1(_036_),
    .C1(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nand2_1 _143_ (.A(_098_),
    .B(_107_),
    .Y(_040_));
 sky130_fd_sc_hd__a31o_1 _144_ (.A1(\bit_idx[2] ),
    .A2(\bit_idx[1] ),
    .A3(\bit_idx[0] ),
    .B1(_040_),
    .X(_041_));
 sky130_fd_sc_hd__or4_1 _145_ (.A(\state[2] ),
    .B(\state[0] ),
    .C(_098_),
    .D(net10),
    .X(_042_));
 sky130_fd_sc_hd__and3_1 _146_ (.A(_039_),
    .B(_041_),
    .C(_042_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _147_ (.A0(\state[0] ),
    .A1(_107_),
    .S(_043_),
    .X(_044_));
 sky130_fd_sc_hd__clkbuf_1 _148_ (.A(_044_),
    .X(_003_));
 sky130_fd_sc_hd__buf_2 _149_ (.A(_039_),
    .X(_045_));
 sky130_fd_sc_hd__and4_1 _150_ (.A(_108_),
    .B(_045_),
    .C(_041_),
    .D(_042_),
    .X(_046_));
 sky130_fd_sc_hd__and4b_1 _151_ (.A_N(_107_),
    .B(_045_),
    .C(_042_),
    .D(_098_),
    .X(_047_));
 sky130_fd_sc_hd__o21ba_1 _152_ (.A1(_098_),
    .A2(_046_),
    .B1_N(_047_),
    .X(_004_));
 sky130_fd_sc_hd__a2bb2o_1 _153_ (.A1_N(_102_),
    .A2_N(_043_),
    .B1(_046_),
    .B2(_098_),
    .X(_005_));
 sky130_fd_sc_hd__a31o_1 _154_ (.A1(\clk_cnt[8] ),
    .A2(\clk_cnt[7] ),
    .A3(_034_),
    .B1(_036_),
    .X(_048_));
 sky130_fd_sc_hd__nor2_1 _155_ (.A(_048_),
    .B(_038_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_2 _156_ (.A(_037_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _157_ (.A0(_049_),
    .A1(_050_),
    .S(\clk_cnt[0] ),
    .X(_051_));
 sky130_fd_sc_hd__clkbuf_1 _158_ (.A(_051_),
    .X(_006_));
 sky130_fd_sc_hd__o21bai_1 _159_ (.A1(\clk_cnt[0] ),
    .A2(_045_),
    .B1_N(_037_),
    .Y(_052_));
 sky130_fd_sc_hd__or3b_1 _160_ (.A(_045_),
    .B(\clk_cnt[1] ),
    .C_N(\clk_cnt[0] ),
    .X(_053_));
 sky130_fd_sc_hd__a21bo_1 _161_ (.A1(net26),
    .A2(_052_),
    .B1_N(_053_),
    .X(_007_));
 sky130_fd_sc_hd__a21o_1 _162_ (.A1(\clk_cnt[1] ),
    .A2(\clk_cnt[0] ),
    .B1(\clk_cnt[2] ),
    .X(_054_));
 sky130_fd_sc_hd__nand3_1 _163_ (.A(\clk_cnt[1] ),
    .B(\clk_cnt[2] ),
    .C(\clk_cnt[0] ),
    .Y(_055_));
 sky130_fd_sc_hd__a32o_1 _164_ (.A1(_049_),
    .A2(_054_),
    .A3(_055_),
    .B1(_050_),
    .B2(net21),
    .X(_008_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(net23),
    .Y(_056_));
 sky130_fd_sc_hd__and4_1 _166_ (.A(\clk_cnt[3] ),
    .B(\clk_cnt[1] ),
    .C(\clk_cnt[2] ),
    .D(\clk_cnt[0] ),
    .X(_057_));
 sky130_fd_sc_hd__o2bb2a_1 _167_ (.A1_N(\clk_cnt[3] ),
    .A2_N(_037_),
    .B1(_045_),
    .B2(_057_),
    .X(_058_));
 sky130_fd_sc_hd__a21oi_1 _168_ (.A1(_056_),
    .A2(_055_),
    .B1(_058_),
    .Y(_009_));
 sky130_fd_sc_hd__and2_1 _169_ (.A(\clk_cnt[4] ),
    .B(_057_),
    .X(_059_));
 sky130_fd_sc_hd__nor2_1 _170_ (.A(_045_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__o21bai_1 _171_ (.A1(_045_),
    .A2(_059_),
    .B1_N(_037_),
    .Y(_061_));
 sky130_fd_sc_hd__a22o_1 _172_ (.A1(_057_),
    .A2(_060_),
    .B1(_061_),
    .B2(net19),
    .X(_010_));
 sky130_fd_sc_hd__or3b_1 _173_ (.A(\clk_cnt[5] ),
    .B(_045_),
    .C_N(_059_),
    .X(_062_));
 sky130_fd_sc_hd__a21bo_1 _174_ (.A1(net34),
    .A2(_061_),
    .B1_N(_062_),
    .X(_011_));
 sky130_fd_sc_hd__a31o_1 _175_ (.A1(\clk_cnt[5] ),
    .A2(\clk_cnt[4] ),
    .A3(_057_),
    .B1(\clk_cnt[6] ),
    .X(_063_));
 sky130_fd_sc_hd__nand3_1 _176_ (.A(\clk_cnt[6] ),
    .B(\clk_cnt[5] ),
    .C(_059_),
    .Y(_064_));
 sky130_fd_sc_hd__a32o_1 _177_ (.A1(_049_),
    .A2(_063_),
    .A3(_064_),
    .B1(_050_),
    .B2(net22),
    .X(_012_));
 sky130_fd_sc_hd__and4_1 _178_ (.A(\clk_cnt[7] ),
    .B(\clk_cnt[6] ),
    .C(\clk_cnt[5] ),
    .D(_059_),
    .X(_065_));
 sky130_fd_sc_hd__o21bai_1 _179_ (.A1(_045_),
    .A2(_065_),
    .B1_N(_037_),
    .Y(_066_));
 sky130_fd_sc_hd__or3_1 _180_ (.A(\clk_cnt[7] ),
    .B(_045_),
    .C(_064_),
    .X(_067_));
 sky130_fd_sc_hd__a21bo_1 _181_ (.A1(net20),
    .A2(_066_),
    .B1_N(_067_),
    .X(_013_));
 sky130_fd_sc_hd__a22o_1 _182_ (.A1(_049_),
    .A2(_065_),
    .B1(_066_),
    .B2(net18),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net24),
    .B(_050_),
    .X(_068_));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(_068_),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _185_ (.A(net32),
    .B(_050_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _186_ (.A(_069_),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net25),
    .B(_050_),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(_070_),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _189_ (.A(net28),
    .B(_050_),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(_071_),
    .X(_018_));
 sky130_fd_sc_hd__and2_1 _191_ (.A(net29),
    .B(_050_),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(_072_),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _193_ (.A(net30),
    .B(_050_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(_073_),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _195_ (.A(net27),
    .B(_050_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(_074_),
    .X(_021_));
 sky130_fd_sc_hd__and3_1 _197_ (.A(_098_),
    .B(_107_),
    .C(_048_),
    .X(_075_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(_098_),
    .Y(_076_));
 sky130_fd_sc_hd__o21ai_1 _199_ (.A1(_076_),
    .A2(_048_),
    .B1(_107_),
    .Y(_077_));
 sky130_fd_sc_hd__mux2_1 _200_ (.A0(_075_),
    .A1(_077_),
    .S(\bit_idx[0] ),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_1 _201_ (.A(_078_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_1 _202_ (.A(\bit_idx[1] ),
    .B(\bit_idx[0] ),
    .Y(_079_));
 sky130_fd_sc_hd__or2_1 _203_ (.A(\bit_idx[1] ),
    .B(\bit_idx[0] ),
    .X(_080_));
 sky130_fd_sc_hd__a32o_1 _204_ (.A1(_079_),
    .A2(_075_),
    .A3(_080_),
    .B1(_077_),
    .B2(net31),
    .X(_023_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(_041_),
    .Y(_081_));
 sky130_fd_sc_hd__o2111a_1 _206_ (.A1(_076_),
    .A2(_048_),
    .B1(_107_),
    .C1(\bit_idx[0] ),
    .D1(\bit_idx[1] ),
    .X(_082_));
 sky130_fd_sc_hd__o22a_1 _207_ (.A1(_081_),
    .A2(_077_),
    .B1(_082_),
    .B2(net17),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _208_ (.A0(net1),
    .A1(net35),
    .S(_100_),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(_083_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _210_ (.A0(net2),
    .A1(net39),
    .S(_100_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(_084_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _212_ (.A0(net3),
    .A1(net41),
    .S(_100_),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_1 _213_ (.A(_085_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _214_ (.A0(net4),
    .A1(net37),
    .S(_100_),
    .X(_086_));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(_086_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _216_ (.A0(net5),
    .A1(net36),
    .S(_100_),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_1 _217_ (.A(_087_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _218_ (.A0(net6),
    .A1(net33),
    .S(_100_),
    .X(_088_));
 sky130_fd_sc_hd__clkbuf_1 _219_ (.A(_088_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _220_ (.A0(net7),
    .A1(net42),
    .S(_100_),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_1 _221_ (.A(_089_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _222_ (.A0(net8),
    .A1(net38),
    .S(_100_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _223_ (.A(_090_),
    .X(_032_));
 sky130_fd_sc_hd__dfrtp_1 _224_ (.CLK(clknet_2_1__leaf_clk),
    .D(_000_),
    .RESET_B(net13),
    .Q(parity_bit));
 sky130_fd_sc_hd__dfstp_1 _225_ (.CLK(clknet_2_1__leaf_clk),
    .D(_001_),
    .SET_B(net15),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_2 _226_ (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .RESET_B(net16),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_4 _227_ (.CLK(clknet_2_3__leaf_clk),
    .D(_003_),
    .RESET_B(net16),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _228_ (.CLK(clknet_2_3__leaf_clk),
    .D(_004_),
    .RESET_B(net16),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _229_ (.CLK(clknet_2_3__leaf_clk),
    .D(_005_),
    .RESET_B(net16),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _230_ (.CLK(clknet_2_2__leaf_clk),
    .D(_006_),
    .RESET_B(net15),
    .Q(\clk_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _231_ (.CLK(clknet_2_2__leaf_clk),
    .D(_007_),
    .RESET_B(net15),
    .Q(\clk_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _232_ (.CLK(clknet_2_2__leaf_clk),
    .D(_008_),
    .RESET_B(net15),
    .Q(\clk_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _233_ (.CLK(clknet_2_2__leaf_clk),
    .D(_009_),
    .RESET_B(net15),
    .Q(\clk_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _234_ (.CLK(clknet_2_2__leaf_clk),
    .D(_010_),
    .RESET_B(net15),
    .Q(\clk_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _235_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .RESET_B(net15),
    .Q(\clk_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _236_ (.CLK(clknet_2_2__leaf_clk),
    .D(_012_),
    .RESET_B(net15),
    .Q(\clk_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _237_ (.CLK(clknet_2_3__leaf_clk),
    .D(_013_),
    .RESET_B(net15),
    .Q(\clk_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _238_ (.CLK(clknet_2_3__leaf_clk),
    .D(_014_),
    .RESET_B(net15),
    .Q(\clk_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _239_ (.CLK(clknet_2_2__leaf_clk),
    .D(_015_),
    .RESET_B(net13),
    .Q(\clk_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _240_ (.CLK(clknet_2_0__leaf_clk),
    .D(_016_),
    .RESET_B(net13),
    .Q(\clk_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _241_ (.CLK(clknet_2_0__leaf_clk),
    .D(_017_),
    .RESET_B(net13),
    .Q(\clk_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _242_ (.CLK(clknet_2_0__leaf_clk),
    .D(_018_),
    .RESET_B(net13),
    .Q(\clk_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _243_ (.CLK(clknet_2_0__leaf_clk),
    .D(_019_),
    .RESET_B(net13),
    .Q(\clk_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _244_ (.CLK(clknet_2_0__leaf_clk),
    .D(_020_),
    .RESET_B(net13),
    .Q(\clk_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _245_ (.CLK(clknet_2_2__leaf_clk),
    .D(_021_),
    .RESET_B(net13),
    .Q(\clk_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_4 _246_ (.CLK(clknet_2_0__leaf_clk),
    .D(_022_),
    .RESET_B(net13),
    .Q(\bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_2 _247_ (.CLK(clknet_2_0__leaf_clk),
    .D(_023_),
    .RESET_B(net13),
    .Q(\bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _248_ (.CLK(clknet_2_1__leaf_clk),
    .D(_024_),
    .RESET_B(net14),
    .Q(\bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _249_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .RESET_B(net14),
    .Q(\data_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _250_ (.CLK(clknet_2_1__leaf_clk),
    .D(_026_),
    .RESET_B(net14),
    .Q(\data_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _251_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .RESET_B(net14),
    .Q(\data_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _252_ (.CLK(clknet_2_1__leaf_clk),
    .D(_028_),
    .RESET_B(net14),
    .Q(\data_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _253_ (.CLK(clknet_2_0__leaf_clk),
    .D(_029_),
    .RESET_B(net14),
    .Q(\data_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _254_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .RESET_B(net14),
    .Q(\data_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _255_ (.CLK(clknet_2_1__leaf_clk),
    .D(_031_),
    .RESET_B(net14),
    .Q(\data_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _256_ (.CLK(clknet_2_1__leaf_clk),
    .D(_032_),
    .RESET_B(net14),
    .Q(\data_reg[7] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(data_in[1]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(data_in[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(data_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(data_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(data_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(data_in[6]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(data_in[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(rst_n),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(tx_start),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(tx_busy));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(tx_out));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net16),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(net9),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\bit_idx[2] ),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\clk_cnt[8] ),
    .X(net18));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\clk_cnt[4] ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\clk_cnt[7] ),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\clk_cnt[2] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\clk_cnt[6] ),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\clk_cnt[3] ),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\clk_cnt[9] ),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\clk_cnt[11] ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\clk_cnt[1] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\clk_cnt[15] ),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\clk_cnt[12] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\clk_cnt[13] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\clk_cnt[14] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\bit_idx[1] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\clk_cnt[10] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\data_reg[5] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\clk_cnt[5] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\data_reg[0] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\data_reg[4] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\data_reg[3] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\data_reg[7] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\data_reg[1] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(parity_bit),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\data_reg[2] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\data_reg[6] ),
    .X(net42));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_293 ();
endmodule
